--same as tb for and gate. reason same no of input and outputs
library ieee;
use ieee.std_logic_1164.all;

entity tb_or_gate is
end entity;

architecture sim of tb_or_gate is
  signal a, b, y : std_logic;
begin
  -- Instantiate the DUT
  uut: entity work.or_gate
    port map (
      a => a,
      b => b,
      y => y
    );

  -- Stimulus process
  process
  begin
    a <= '0'; b <= '0'; wait for 100 fs;
    a <= '0'; b <= '1'; wait for 100 fs;
    a <= '1'; b <= '0'; wait for 100 fs;
    a <= '1'; b <= '1'; wait for 100 fs;
    wait;  -- stop simulation
  end process;
end architecture;
